library verilog;
use verilog.vl_types.all;
entity proc2 is
    generic(
        T0              : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        T1              : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi1);
        T2              : vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi0);
        T3              : vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi1);
        T4              : vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi0);
        T5              : vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi1);
        b               : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        beq             : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi1);
        bne             : vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi0);
        mv              : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        mvt_b           : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi1);
        add             : vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi0);
        sub             : vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi1);
        ld              : vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi0);
        st              : vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi1);
        \And\           : vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi0);
        shift_rot       : vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi1);
        R0              : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        R1              : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi1);
        R2              : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi1, Hi0);
        R3              : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi1, Hi1);
        R4              : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi0);
        R5              : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi1);
        R6              : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi1, Hi0);
        PC              : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi1, Hi1);
        G               : vl_logic_vector(0 to 3) := (Hi1, Hi0, Hi0, Hi0);
        IR8_IR8_0       : vl_logic_vector(0 to 3) := (Hi1, Hi0, Hi0, Hi1);
        IR7_0_0         : vl_logic_vector(0 to 3) := (Hi1, Hi0, Hi1, Hi0);
        data            : vl_logic_vector(0 to 3) := (Hi1, Hi0, Hi1, Hi1)
    );
    port(
        Resetn          : in     vl_logic;
        Clock           : in     vl_logic;
        Run             : in     vl_logic;
        Done            : out    vl_logic;
        \_r0\           : out    vl_logic_vector(15 downto 0);
        \_r1\           : out    vl_logic_vector(15 downto 0);
        \_r2\           : out    vl_logic_vector(15 downto 0);
        \_r3\           : out    vl_logic_vector(15 downto 0);
        \_r4\           : out    vl_logic_vector(15 downto 0);
        \_pc\           : out    vl_logic_vector(15 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of T0 : constant is 1;
    attribute mti_svvh_generic_type of T1 : constant is 1;
    attribute mti_svvh_generic_type of T2 : constant is 1;
    attribute mti_svvh_generic_type of T3 : constant is 1;
    attribute mti_svvh_generic_type of T4 : constant is 1;
    attribute mti_svvh_generic_type of T5 : constant is 1;
    attribute mti_svvh_generic_type of b : constant is 1;
    attribute mti_svvh_generic_type of beq : constant is 1;
    attribute mti_svvh_generic_type of bne : constant is 1;
    attribute mti_svvh_generic_type of mv : constant is 1;
    attribute mti_svvh_generic_type of mvt_b : constant is 1;
    attribute mti_svvh_generic_type of add : constant is 1;
    attribute mti_svvh_generic_type of sub : constant is 1;
    attribute mti_svvh_generic_type of ld : constant is 1;
    attribute mti_svvh_generic_type of st : constant is 1;
    attribute mti_svvh_generic_type of \And\ : constant is 1;
    attribute mti_svvh_generic_type of shift_rot : constant is 1;
    attribute mti_svvh_generic_type of R0 : constant is 1;
    attribute mti_svvh_generic_type of R1 : constant is 1;
    attribute mti_svvh_generic_type of R2 : constant is 1;
    attribute mti_svvh_generic_type of R3 : constant is 1;
    attribute mti_svvh_generic_type of R4 : constant is 1;
    attribute mti_svvh_generic_type of R5 : constant is 1;
    attribute mti_svvh_generic_type of R6 : constant is 1;
    attribute mti_svvh_generic_type of PC : constant is 1;
    attribute mti_svvh_generic_type of G : constant is 1;
    attribute mti_svvh_generic_type of IR8_IR8_0 : constant is 1;
    attribute mti_svvh_generic_type of IR7_0_0 : constant is 1;
    attribute mti_svvh_generic_type of data : constant is 1;
end proc2;
